module Macro_Tb ();
  reg Clk,Rst,WE;
  reg [63:0]BL,BLB;
  reg Addr;
  reg [127:0]WL;
  reg [127:0]In_B;
  reg wb;
  wire [63:0]DOut;
  
  
 initial
  begin
    Clk=1'b1;
    Rst=1'b1;
    WE=1'b1;
    BL=64'b1111111111111111111111111111111111111111111111111111111111111111;
   BLB=64'b0000000000000000000000000000000000000000000000000000000000000000;
   Addr=1'b1;
   WL=128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
 In_B=128'b10000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000;
 wb=1'b1;
 
 #500
 
 Rst=1'b0;
 
 
   
    
   
#500
$finish; 


end


   initial
   begin
     
     
     
   
     $dumpfile("Macro_SXAFA.vcd");
     $dumpvars;
     
   end 
   
   
   Macro M0 (Clk,Rst,WE,BL,BLB,Addr,WL,In_B,wb,DOut);
   
 endmodule